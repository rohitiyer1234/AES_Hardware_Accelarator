module RoundKey_mem(
    input clk, reset
);
endmodule